`include "packet_if.svi"

module hw_top;

packet_if vif();

endmodule

