`ifndef __PACKET_DEFINE_SV__
`define __PACKET_DEFINE_SV__

`include "packet.sv"

typedef mailbox #(packet) packet_tran_mbox;

`endif

